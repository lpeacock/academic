module data_flow(
    input [7:0] x_in,
    output [7:0] y_out
    );
endmodule
